`define PRECISION 8
`define CSIZE 9
`define CROW 3